`include "../src/parameter.v"

module LDED( // Largest and Duplicate Element Detector
    input rst,
    input clk_mn,
    input [`ELEMENT_NUM-1:0] FO_mj_reg,
    input mode,
    input mj_level,
    output SM_valid,
    output reg TR_empty, // reg, output to mj
    output reg [`LOG2_ELEMENT_NUM-1:0] LE_Addr // wire
);

// assume clk_mj > 4 * clk_mn ??

reg mn_level_sync[0:2];
wire mn_pulse = mn_level_sync[1] ^ mn_level_sync[2]; // XOR

reg [`ELEMENT_NUM-1:0] Temp_Reg;
reg [`ELEMENT_NUM-1:0] TR_nxt;

// wait for mn_pulse, which means FO_mj_reg is stable
wire [`ELEMENT_NUM-1:0] TR_comb = (mn_pulse)? FO_mj_reg: Temp_Reg;

wire one_one = (|TR_comb) && (TR_comb == (TR_comb & -TR_comb));
assign SM_valid = |TR_comb;

// minor clock domain
always@(posedge clk_mn) begin
    if(rst) begin
        Temp_Reg <= 0;
        TR_empty <= 1;
    end
    else if(mode) begin // Sorting output mode
        Temp_Reg <= TR_nxt;

        // if there is one left in TR, then next cycle set empty=1
        TR_empty <= (!SM_valid || one_one)? 1: 0;
    end
end

always@(posedge clk_mn) begin
    mn_level_sync[0] <= mj_level; // mn_level_sync[0] may be metastable
    mn_level_sync[1] <= mn_level_sync[0]; // mn_level_sync[1] won't be metastable
    mn_level_sync[2] <= mn_level_sync[1];
end

always@(*) begin
    // assume ELEMENT_NUM = 16
    // 16 ELEMENT DECODER
    TR_nxt = TR_comb;
    casez(TR_comb)
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1: begin LE_Addr = 0;	TR_nxt[0]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10: begin LE_Addr = 1;	TR_nxt[1]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100: begin LE_Addr = 2;	TR_nxt[2]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000: begin LE_Addr = 3;	TR_nxt[3]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000: begin LE_Addr = 4;	TR_nxt[4]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000: begin LE_Addr = 5;	TR_nxt[5]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000: begin LE_Addr = 6;	TR_nxt[6]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000: begin LE_Addr = 7;	TR_nxt[7]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000: begin LE_Addr = 8;	TR_nxt[8]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000: begin LE_Addr = 9;	TR_nxt[9]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000: begin LE_Addr = 10;	TR_nxt[10]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000: begin LE_Addr = 11;	TR_nxt[11]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000: begin LE_Addr = 12;	TR_nxt[12]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000: begin LE_Addr = 13;	TR_nxt[13]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000: begin LE_Addr = 14;	TR_nxt[14]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000: begin LE_Addr = 15;	TR_nxt[15]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000: begin LE_Addr = 16;	TR_nxt[16]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000: begin LE_Addr = 17;	TR_nxt[17]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000: begin LE_Addr = 18;	TR_nxt[18]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000: begin LE_Addr = 19;	TR_nxt[19]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000: begin LE_Addr = 20;	TR_nxt[20]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000: begin LE_Addr = 21;	TR_nxt[21]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000: begin LE_Addr = 22;	TR_nxt[22]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000: begin LE_Addr = 23;	TR_nxt[23]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000: begin LE_Addr = 24;	TR_nxt[24]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000: begin LE_Addr = 25;	TR_nxt[25]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000: begin LE_Addr = 26;	TR_nxt[26]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 27;	TR_nxt[27]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 28;	TR_nxt[28]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 29;	TR_nxt[29]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 30;	TR_nxt[30]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 31;	TR_nxt[31]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 32;	TR_nxt[32]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 33;	TR_nxt[33]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 34;	TR_nxt[34]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 35;	TR_nxt[35]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 36;	TR_nxt[36]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 37;	TR_nxt[37]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 38;	TR_nxt[38]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 39;	TR_nxt[39]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 40;	TR_nxt[40]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 41;	TR_nxt[41]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 42;	TR_nxt[42]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 43;	TR_nxt[43]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 44;	TR_nxt[44]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 45;	TR_nxt[45]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 46;	TR_nxt[46]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 47;	TR_nxt[47]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 48;	TR_nxt[48]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 49;	TR_nxt[49]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 50;	TR_nxt[50]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 51;	TR_nxt[51]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 52;	TR_nxt[52]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 53;	TR_nxt[53]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 54;	TR_nxt[54]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 55;	TR_nxt[55]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 56;	TR_nxt[56]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 57;	TR_nxt[57]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 58;	TR_nxt[58]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 59;	TR_nxt[59]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 60;	TR_nxt[60]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 61;	TR_nxt[61]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 62;	TR_nxt[62]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 63;	TR_nxt[63]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 64;	TR_nxt[64]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 65;	TR_nxt[65]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 66;	TR_nxt[66]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 67;	TR_nxt[67]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 68;	TR_nxt[68]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 69;	TR_nxt[69]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 70;	TR_nxt[70]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 71;	TR_nxt[71]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 72;	TR_nxt[72]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 73;	TR_nxt[73]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 74;	TR_nxt[74]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 75;	TR_nxt[75]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 76;	TR_nxt[76]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 77;	TR_nxt[77]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 78;	TR_nxt[78]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 79;	TR_nxt[79]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 80;	TR_nxt[80]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 81;	TR_nxt[81]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 82;	TR_nxt[82]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 83;	TR_nxt[83]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 84;	TR_nxt[84]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 85;	TR_nxt[85]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 86;	TR_nxt[86]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 87;	TR_nxt[87]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 88;	TR_nxt[88]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 89;	TR_nxt[89]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 90;	TR_nxt[90]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 91;	TR_nxt[91]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 92;	TR_nxt[92]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 93;	TR_nxt[93]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 94;	TR_nxt[94]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 95;	TR_nxt[95]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 96;	TR_nxt[96]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 97;	TR_nxt[97]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 98;	TR_nxt[98]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 99;	TR_nxt[99]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 100;	TR_nxt[100]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 101;	TR_nxt[101]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 102;	TR_nxt[102]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 103;	TR_nxt[103]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 104;	TR_nxt[104]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 105;	TR_nxt[105]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 106;	TR_nxt[106]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 107;	TR_nxt[107]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 108;	TR_nxt[108]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 109;	TR_nxt[109]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 110;	TR_nxt[110]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 111;	TR_nxt[111]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 112;	TR_nxt[112]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 113;	TR_nxt[113]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 114;	TR_nxt[114]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 115;	TR_nxt[115]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 116;	TR_nxt[116]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 117;	TR_nxt[117]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 118;	TR_nxt[118]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 119;	TR_nxt[119]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 120;	TR_nxt[120]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 121;	TR_nxt[121]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 122;	TR_nxt[122]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 123;	TR_nxt[123]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 124;	TR_nxt[124]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 125;	TR_nxt[125]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 126;	TR_nxt[126]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 127;	TR_nxt[127]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 128;	TR_nxt[128]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 129;	TR_nxt[129]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 130;	TR_nxt[130]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 131;	TR_nxt[131]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 132;	TR_nxt[132]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 133;	TR_nxt[133]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 134;	TR_nxt[134]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 135;	TR_nxt[135]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 136;	TR_nxt[136]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 137;	TR_nxt[137]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 138;	TR_nxt[138]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 139;	TR_nxt[139]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 140;	TR_nxt[140]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 141;	TR_nxt[141]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 142;	TR_nxt[142]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 143;	TR_nxt[143]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 144;	TR_nxt[144]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 145;	TR_nxt[145]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 146;	TR_nxt[146]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 147;	TR_nxt[147]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 148;	TR_nxt[148]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 149;	TR_nxt[149]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 150;	TR_nxt[150]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 151;	TR_nxt[151]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 152;	TR_nxt[152]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 153;	TR_nxt[153]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 154;	TR_nxt[154]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 155;	TR_nxt[155]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 156;	TR_nxt[156]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 157;	TR_nxt[157]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 158;	TR_nxt[158]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 159;	TR_nxt[159]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 160;	TR_nxt[160]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 161;	TR_nxt[161]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 162;	TR_nxt[162]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 163;	TR_nxt[163]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 164;	TR_nxt[164]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 165;	TR_nxt[165]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 166;	TR_nxt[166]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 167;	TR_nxt[167]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 168;	TR_nxt[168]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 169;	TR_nxt[169]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 170;	TR_nxt[170]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 171;	TR_nxt[171]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 172;	TR_nxt[172]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 173;	TR_nxt[173]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 174;	TR_nxt[174]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 175;	TR_nxt[175]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 176;	TR_nxt[176]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 177;	TR_nxt[177]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 178;	TR_nxt[178]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 179;	TR_nxt[179]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 180;	TR_nxt[180]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 181;	TR_nxt[181]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 182;	TR_nxt[182]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 183;	TR_nxt[183]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 184;	TR_nxt[184]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 185;	TR_nxt[185]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 186;	TR_nxt[186]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 187;	TR_nxt[187]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 188;	TR_nxt[188]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 189;	TR_nxt[189]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 190;	TR_nxt[190]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 191;	TR_nxt[191]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 192;	TR_nxt[192]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 193;	TR_nxt[193]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 194;	TR_nxt[194]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 195;	TR_nxt[195]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 196;	TR_nxt[196]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 197;	TR_nxt[197]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 198;	TR_nxt[198]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 199;	TR_nxt[199]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 200;	TR_nxt[200]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 201;	TR_nxt[201]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 202;	TR_nxt[202]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 203;	TR_nxt[203]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 204;	TR_nxt[204]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 205;	TR_nxt[205]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 206;	TR_nxt[206]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 207;	TR_nxt[207]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 208;	TR_nxt[208]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 209;	TR_nxt[209]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 210;	TR_nxt[210]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 211;	TR_nxt[211]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 212;	TR_nxt[212]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 213;	TR_nxt[213]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 214;	TR_nxt[214]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 215;	TR_nxt[215]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 216;	TR_nxt[216]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 217;	TR_nxt[217]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 218;	TR_nxt[218]	= 0; end
        256'b????_????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 219;	TR_nxt[219]	= 0; end
        256'b????_????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 220;	TR_nxt[220]	= 0; end
        256'b????_????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 221;	TR_nxt[221]	= 0; end
        256'b????_????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 222;	TR_nxt[222]	= 0; end
        256'b????_????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 223;	TR_nxt[223]	= 0; end
        256'b????_????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 224;	TR_nxt[224]	= 0; end
        256'b????_????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 225;	TR_nxt[225]	= 0; end
        256'b????_????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 226;	TR_nxt[226]	= 0; end
        256'b????_????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 227;	TR_nxt[227]	= 0; end
        256'b????_????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 228;	TR_nxt[228]	= 0; end
        256'b????_????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 229;	TR_nxt[229]	= 0; end
        256'b????_????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 230;	TR_nxt[230]	= 0; end
        256'b????_????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 231;	TR_nxt[231]	= 0; end
        256'b????_????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 232;	TR_nxt[232]	= 0; end
        256'b????_????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 233;	TR_nxt[233]	= 0; end
        256'b????_????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 234;	TR_nxt[234]	= 0; end
        256'b????_????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 235;	TR_nxt[235]	= 0; end
        256'b????_????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 236;	TR_nxt[236]	= 0; end
        256'b????_????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 237;	TR_nxt[237]	= 0; end
        256'b????_????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 238;	TR_nxt[238]	= 0; end
        256'b????_????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 239;	TR_nxt[239]	= 0; end
        256'b????_????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 240;	TR_nxt[240]	= 0; end
        256'b????_????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 241;	TR_nxt[241]	= 0; end
        256'b????_????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 242;	TR_nxt[242]	= 0; end
        256'b????_????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 243;	TR_nxt[243]	= 0; end
        256'b????_????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 244;	TR_nxt[244]	= 0; end
        256'b????_????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 245;	TR_nxt[245]	= 0; end
        256'b????_????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 246;	TR_nxt[246]	= 0; end
        256'b????_????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 247;	TR_nxt[247]	= 0; end
        256'b????_???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 248;	TR_nxt[248]	= 0; end
        256'b????_??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 249;	TR_nxt[249]	= 0; end
        256'b????_?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 250;	TR_nxt[250]	= 0; end
        256'b????_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 251;	TR_nxt[251]	= 0; end
        256'b???1_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 252;	TR_nxt[252]	= 0; end
        256'b??10_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 253;	TR_nxt[253]	= 0; end
        256'b?100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 254;	TR_nxt[254]	= 0; end
        256'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: begin LE_Addr = 255;	TR_nxt[255]	= 0; end
        default: begin LE_Addr = 0;	TR_nxt	= 0; end
    endcase

end

endmodule